module Serial_Twos_Comp (output y, input [7: 0] data, input load, shift_control, Clock, reset_b);
